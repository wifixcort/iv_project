//4 bit OR module
module OR ( input [3:0] a, b, output [3:0] or_ );
   assign or_ = a|b;
endmodule // OR

