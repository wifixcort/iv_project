//4 bit XOR module 
module XOR ( input [3:0] a, output y );
   assign y = ^a;
endmodule
