//4 bit AND module 
module AND ( input [3:0] a, b, output [3:0] and_ );
   assign and_ = a&b;
endmodule


   
