//4 bit OR module
module OR ( input [3:0] a, output y );
   assing y = |(a);
endmodule
