//4 bit AND module 
module AND ( input [3:0]a, output y );
   assign y = &(a);
endmodule


   
