//4 bit AND module 
module AND ( input a, output y );
//   assing y = &(a);
   assing y = a;   
endmodule


   
