//4 bit OR module
module OR ( input [3:0] a, output or_ );
   assign or_ = |a;
endmodule
