//4 bit AND module 
module AND ( input [3:0]a, output and_ );
   assign and_ = &(a);
endmodule


   
