//4 bit XOR module 
module XOR ( input [3:0] a, b, output [3:0] xor_ );
   assign xor_ = a^b;
endmodule
